`include "common.sv"
`include "interface.sv"
`include "transaction.sv"
`include "alu_gen.sv"
`include "alu_bfm.sv"
`include "alu_mon.sv"
`include "alu_cov.sv"
`include "alu_agent.sv"
`include "alu_sbd.sv"
`include "alu_env.sv"
`include "module_top.sv"
