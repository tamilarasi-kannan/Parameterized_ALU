interface alu_int();
  bit [n-1:0]a,b;
  bit [n:0]result;
  bit [2:0] opcode;
endinterface
