mailbox gen2bfm=new();
mailbox mon2cov=new();
mailbox mon2sbd=new();
parameter n=4;
static int num_matches;  
static int num_miss_matches;
static int  count=3 ;
